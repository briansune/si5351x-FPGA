// =====================================================================
//  ____         _                 ____                      
// | __ )  _ __ (_)  __ _  _ __   / ___|  _   _  _ __    ___ 
// |  _ \ | '__|| | / _` || '_ \  \___ \ | | | || '_ \  / _ \
// | |_) || |   | || (_| || | | |  ___) || |_| || | | ||  __/
// |____/ |_|   |_| \__,_||_| |_| |____/  \__,_||_| |_| \___|
// 
// =====================================================================

// module si5351_iic #(
	// parameter system_clk_freq = 100000,
	// parameter [0 : 0] si5351_a0 = 1'b0
// )(
	
	// input			sys_clk,
	// input 			sys_nrst,
	
	// output			ready,
	
	// output			scl,
	// inout			sda
// );


`timescale 1ns / 1ps




`pragma protect begin_protected
`pragma protect version=2
`pragma protect encrypt_agent="ipecrypt"
`pragma protect author="Brian Sune"
`pragma protect author_info="briansune@gmail.com"
`pragma protect data_method="aes128-cbc"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption="true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2020_08"
`pragma protect key_method="rsa"
`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control xilinx_schematic_visibility="false"
`pragma protect control decryption="true"
`pragma protect key_block
A8kudsP17miNhbBYDq5PqEQ6jetO9KN284bdRnR3UhrzpCZkf5uYn4K34gsVlgHb
o5kFJo0TCKnES49u9/AGU/5Bplhb9WreFsrKqbiF0uzoSkzK111+MYkDuuW6ENfa
Q/KcezeAOtJfpaOILE/wpXuO9QL2HgKmYDaIG1yEqMoNQNykoZ7zyiwpi+KMU8aI
jn25QAv4T1qSxgadKESEY5Cl8n0zCKGzPe2vNJi5Qmtkq/HRe1n/dpS29aTZoTXL
lN5e64jnDloVFcB/F4zSL0GHS6FcUNh9R8AhO38KTD5Afnl6MBUfpdMrT8oytUIM
+KldDkgv7oPjbeN+UDJYGA==
`pragma protect end_toolblock="YtASTThKSZSBDafNfI6uTNdiQidGM4fhMcqoS8b0spk="
`pragma protect data_block
LM615/lhrYQ/hSiS2nI/R4a1JXu+iVFbe1sGUBDuks4bg+5km/JJUH/O7CPje4c8
m5tmDo7MSjYQSzHI9u904z2zXVsK1dz5GuaClsOAacq4WfEYVpsyZbOm/DlFaPcU
Lu/laP8f7MD6vf2+c635Wa8lpsXfhzuIBncl3Kttn9jObpXUNvkVPqiCD4Zo6qNY
zXQwJlPZsBZXOQLhxzNaJsXx+rDCiNHLaZhFlLFZUXNDzeYGYc3mEOhUUGFYI3oz
6izx5vno/LgyhrNEL+xOoITkdUoitQd2nFIgyR7PlcHEL9E1LSHvqXno+mdHraUc
/SPzAGmNLm8LYZlnv7NsdGyIYWCzaiI3fylz+hmA95bIEqtq0OrRMnCBQRez6LUm
pn3+PuEvBTpECDByV1R8uGLPUmKFdHAV2ZPR1/IkdntQfW0Ellc+V1F/a30SXTt9
bK7GNIxzWe2HbVS5rlX5PzHB74J58xf1liyD1a1+Xgc0EKzZRLQkpT5nd07mZSAA
6YZeLlpAByLtoZxhtbQ9n3Tk1KCNLt5djAaosRJtYdp8sIXcBnIEJ1uPyCU1ga1S
UVW5cwC+Enor4P4Et+nXwevkYNK+lzV3K+jsgWNIBcogVlXht0XpzzYXhp14Scz0
3O7yE04dTfoNbiggT0hGXlvO5zizzN96mbHZHnuVEUGZYhkM09rb6VYqrEo/oooL
ESge6bBopA+ilzMOW35iuUWqIkqNvwOhqFlBLsYWa61zQRjMvI/1Q03FGLflHpT0
v/D+Y1CX7JwTyO1nNbYTjbXVA9LRyl9ALlujKuD9eL+eIaLad8D5rT7fpRPD4WIa
AVd3Iug9PD3uzkmpJR2vXzdvDgbdMaDLXHHN6dUe3LpuXYBlKnDKGM1AIhe8kqmz
GHevp0y1/8SXSpSoZcibkCp1L0/l8Nojj6nRT5EVp2R1YPterogm/j42DK1ur0YT
WiLMnhcbYscZ+cqiXZ/ZKA7PUM7sHJNrYSxPj2tOO+TBU8NfIQ2q5BENZynbUftl
EnbrQIHG87Jf22rJoCvk1UPKgJE+tBZrItScEUlASHvCSNZDSjPYR9WgvKc/RSDM
uulAP44UbIJ0pQcq/DZH/DvPH2hg/EgKDkBLmqAoFdeHtNw5HwwpLZpu4/X3YXkt
D/QC22lQaAhoDchKsyN95dEvA8ra7GDOjhbdr2FCLjjC7FymUUFvFAxWY2Q9JEpy
8vjlvizBDxLj2c2qqIbB0NXSRQq4WS98BwwG7pAa3WiNnr45AeevGm4tXDNvWnq2
TzrJUK9VabqgIii+fOjscamtzmwVtxz19Sm8v2sl5KlNOXGbJlTg3KU+gE1eKIcy
Xub26OnUR9HVuwwvW7+0bhFzutByveEZF8q/pYIWd+fjtQc6vkj/Y7RnfL+ypjgu
MO3yB6l+lTJKJcvhdDD4PghgjAPZP3myyDb6bFICAgaYp0TRn85TpSDlR8KC3fvO
mwXHOIapfJdiCe2AjtWqoazQ1+BqA0zNGrbT/oM0A/h489zIJgI+Pk/yivAhstaK
EMzQ+ZiOcntS6XYAC/7CFO+dzz7HFysK9i3yI0UyGvrHy5b1V9SeVZDdVJx+kLA7
DilBujjk1DsJmi/tRSv9B6P/e50xvlD6ikuu9GzhMs3kyR0L0NJYhcej7q+9VrXg
/VUMsS8J6cP86z4shaqQprp/yhe3EhTEsGohrZI3fS2kiRaBQeY0oMHcgb4ozhic
FT6CiucMl916U/xvTZGGVZbZPMr1x2TltQIH4oeYyGvir7JTzRRFW2Stqp9B+eDv
Je2/lHMBg0Mo5fBaXpUNRJLkXAhivu1ss2c8ZWzww7ySVsQxEn2od0IRBWxOIZRI
GER5641xt3EVFPky3sWRNYVfHgu00N0xpJt1T5DQIhkNopRx1IU+dILpPWZYjVje
B2pyUj26+JkUxmSpQeSI8zwrUsVUpAex97asQ6xlXIdH+bJdiRQ6oL9eHXW9izIx
yf47QGW7pYv2x1mDQCQY+utUmlWj5YBUqisI2iNAZmH9FyqrCLSqylRlr8ldcs2t
oEwJvxiCiCl7RyBznmUhreUNLdGDvS0VeI59BOAqGNes2uEYh9J1EjkILDe21p67
YTcF7SRU+iGo1akS+og2doF0zIX6562aj9GqRjSdy853DuL3E26Idn66X1NohsYM
55iCUMaNd7ieagAoDrjMqN9b6nqHHjn90zIEbZpoCrYE03a9qrCp5LYkAvKL2KMW
ks8vjiGsH7DMaILMCh36NG+Ig/EVcz1HklHsc2iT5gV0I+89sa0sUtJlIgHAO+ol
bUny2KkUxHesEQjpT9ZePNlTlrW9Wp/mEb2QywNQlmNRozQWxTyaPf+4Ga4Na0Hw
kYpHlxVIfqPcVhe7yrZ/1Y9ElyKUzkHd6kTKhd94mdMaI0Lhm1gg32Q1qNiDouTi
T8ka6b6IetcMkquE21RvHDQQVmAQ6L7dwfAp2wFL5h+HgovuUkU0SmRCzXQW0bkF
jdks1XiNmxXgZWEzlY1YYflTJ3tGrCR9H7ujZMB6ir6nbnLPNjzxg13NSF20qfMz
CiGjV6LcwxAU8waeYeGgRSfzHBzOy4gbuzgrt6lWbCGK8AVvNDTEh0juh7yZvoUl
PVPQ3jQXBsL3ITkZfJswE7ma+fx+O1qZs6DHlVQEnqbHoc/0OcuXk5Ew8+9oQdIB
O3xgty4p2npLKErROlvPwG8iu9n+7MyLGfzxk4tZc+DEZj9Y0eAYtlCFJa7j5sK+
PGnLn8AsDTYb4aPJvbQBtpw0/9drAH/1eL/qe+lqqq5arbqDE20mlaT2ddFeUjR9
O30Zi1Bf20pznuj8v+NkOWvhNb/T5/CkyU6doCR5vp8xp94NB1qubYev5AskixRi
hv1qIxsTyhV6s1Ay6oWIt0sBYFTwOKNVCVLzSJ5a6bcsotuNshNetCL8rzDCxulb
zqhx03DYvyfzNgi0mKMAJHrxmPkxEGa2OCms2qyyIC/ba0GeJl/xi1+ev4Unpp0D
bxVYUPkHUHhnlR9FxuTHR2tTSqA/cJNYCEpSrMSm+MB1Z5Vj6oe46to66Z5hrXtP
hlYK6HDcHllThKCh15e9qWb73DAmsRJfLKdGCylOtKPbJ/kWvLQ4+7bm/vVDYf0H
8fKy6lLHe3bkIjq0avClAtGM9VCMqzGCIt0+daniDJttSl7WXesSfbSfVwP9yOL+
60w//lPQi/MniYWHNsnQHwhxi1+5s+p/1JFVrBxDWABfBNlbne7X2J/Bw3+2H6dM
0W7u7jkZxzIcaZueAcYerFc3GoNh+LNIzQaHU0v5GSiQplVT1PVsjceduF0O1w2j
frn+k/rGlQ52dvcyqs8hidxLvtixDPhCwjXOOZ8IPbNlpqx8b3hqwVzSch2JuHtM
7E1kOEPOmlmg03EkqulbTiaEGDmcyvv2+ryi2OkSfa9H/6v/JzFBRj1ypGJQyVoC
L/xE0rH27/Y5IoiB6y3SjnAkx8JDvSELd3BNab5jEpelDcTNYIEEx8Bg7dylCgA3
coa991H37XsMbEl9grOIbwQZLc+4vEy2sR6B/yO3CqRwEB5IdDb6jPfFvXs6n8/W
rdrD03j5ulp4DXmzqC7jQ6Mdv/Hzu9/D8f6pnA4pPe8xVCXEvL+GJj7TWyMB5B4t
5cc8au/XHVZL3XQnj0oyd7DQCjkuAqbgJppqAMV2GJ5EKNozrfmxxzYm3TF3Ye3E
2fPTzJ0MZTMjBM34Bo+dsKfrl5X2pMz+fBNOQKq8PauHbN8iKqZ4mdmvmyWICe2W
O3oFETGdHiftf14KvtKv2jx/+jWX3PRdYFoL+tXri3WvKYuuljnzSPOyxbTjG6BS
deG0fk9nWKhLCSdRH0ZsmRe4xxXFdRf/TOvcVTZ5uiGcXv3aFtqKHp28vJ/D/7Qm
Tmn1sLPIr4/Vqfj94NtNx/tIbupFM/nb0t1NNn9tpQFvIu6SePFxg0LEgusOaBJh
WLtpQTnfS2JsgxH5rJdNTQl7XWV/K0A8wjLOv//y1X+4I/i/mEspNJ5TbUV//Tpt
2YIYXbNjaOkKIMrNgI3n4wl2WdpoCMrg21X+CEdSohcGlApcbFr/o8Yh6Lg7T2IV
J4st5IB9w8NGxm+DosLngQUuYqbm1bgxC4xhKwNgkXpkQ13ODmd8njkFwG2mjcPO
7HZNTAYAVgcX9LlIhej3tO9k3d4MCOzi852lgfs7OvIyXG/dgQ+D0BvWs4ecy63w
8v2IbMhED3UlXdJefzcU229KAItTG5d4wvO2etlp+cUsPrQSej8iWM08bmxUh1Jt
WCjhKDGV1WRfNCh0+j2I+OGINzgLnr3Aspdhw3/eknCHXfWDnKf5SSGtHdK3M0IR
+Bfl5Q4EEHoiftOwF+YJkr/QNRDgJDAS9gnc4Vbl8nlXVcSBqENIInYm66zD3ukb
P0HBh5k3LDVJGNjwloIUgh/esZF2HxufbRrsHO6ZbWl4zKrEBAB8nFno8zc+GL0y
Pp+SJoUtNRAWV9qMI69NMsLE/TC7F7EhrlWAcsFz1bETOdOSLv60ipryj2Aro1zD
0kl9e/eETr+tJnMTVzUY2FxFgqI9+fQKZlr+ibWH409+E8X1ztvu+zVDMvG3qH83
rDVhsMEupLHjJ8wQ4bk3p36AoT8YXt5beuP8/2a0XLtRpA9XeVl2pw1lnZol082x
Nd9xr65CXVSKPkC3nRhtkqbX4OW403SUTiFhQC+mhLD9zE8EfNlRby3OxkFY1jDU
yum6tLKeF9TGyg4fmiz9FXyeITnjEh2OmbynM7RWeE1bFRaVospkOYeGeCvgpqgq
HMLK9NS2jyYG/EDFYQ76hR0mPAIkjfYz5dq1Zp6u7ZIQUOzyzOvjXBnvvvcicUhQ
G4iszApDU+PdQZiF6h2ywEVBVla5nA6B5l7ApxmcJeCdRa00OCmuba0kuQfHn/OT
g2gkqO1DaMLkASoc/YwwUD3aQ44VwmRwWGS41kXxaliO0aUz2+iq6GBGdr9EPZVr
dNBLooNfaoqhW14ATtczUgN+0iQtbuHL/TXw1R+HQc8zHD4p8VzWDvcI3Rtb16vR
YbimyH6+tpX7+bfQKx69mJks6JPySlmVl/kEXbg9s/tQiD2xL3kR22mOm5qb1B2J
vJRRd+RGyVLVvoyIbJN522KSjOs/W9P19uBgosEDErHOj5i0MXrdVCEtuFLZX2Ge
zttdQnwSM+T6Y04VEZKefcWRbNXfVn6aC1YlFLhf0XqGW5P8eY6O0EGvl2JD3teG
jyyOMl/tpoBHtEh2uJS2PsBE6KIcGYY+wc0tBYsEzZ8P8W2dBNPqawIg05RhfFSs
lExgbnwg8o4TMnlZNCmMPMytrcpi6Yo76tqNW6fy/ocvChG7j1CBVFGavv9L9ImL
LwkRBxi6z3TnzgHNVvdQeN+ZbDjSSICU2gi9J/KImYKjpdcSM8yC8VlFfTIr2zPh
w7C/wtPc7IEHz8NmFNtO7C9hHTJ6uX8S7+TWNuzBB7GxxwbvYdZGMV+J/XxMSGbo
JqNqStCUaqfMzztDJjo8Gu8ftXp9eHWqReWFK/J4YK8eAT/OIFhGwhh3gDDTs4+2
sIqPOlkqL92g69uIf7ZiqZ4NJjY6hG1Awx/FWWtjfgOXIlQBZj2ehwa3ghZE3a0Q
wIA7fuM0doXz3V8sbZe6y582lfCR4QnH63wRoWigeca9R6BrDgj6vIzLXylTrw2/
yOWa3pxDc0I+kcI0/JS+ysNnAuWMEdZrKw2hej1cPYJeRuUWlT0QSeOM2F1Ys4OA
i3hCxE6x/YOSJNPLHXVCPS6c9LKTQ8oDcE798kBnkei3Y+axpmmgHZhfVf9Z5e41
ZLUsjc9zSxiZFoGUiBt17Kh9g0C/rB0CKyue1mZmXp4J0D0CHwiyGMc9AUYRrb7c
bXDxhWID1nWGqL9xFjgY9HbIjcjJ7vCHbuaGyawJ1AOCeFzFhka05A7bTzK/VKiM
bOvv5nqd+qi78Abn+PrJinxqFwWB42tvUJgA6NY8YCgbfMOhUB5qFL0MyarnqDHG
QWKMYxQTAWqQ4N/J4PEBaSydP06NRPLYWueox5lLLcbAbgFEW2hbD6lsyxB92Znl
4tDdSnXCOBlhBXl+VIfOgqjxrRf/8E74dH4IB0NuDP1oqLdWg/NKJn/GP4gwI6JX
BjyggZNE5jpGZr/bFiMK6yFfgEM6Qfk+90zzwiCG4elrgLtLtZoXIzf3hO5ip4FG
az3svQKhQgHQv+kYLOJEQk45RO5W1hn5ZNXVecbqCqReZqBVSFZiP/+g6l0pmHDp
pzovVfvBXMcfbPIpCp+yRX5AJAYaKKS9kJL7kkUXU15IDQdB4YH5aK5rWoHDidh/
x4Hx+SAb/aD4hUUgzWRpNMZ2/rUKVQeDnBix9j3g6U5hpVzRbUkv2Z23iPrmAVoC
ZPgZMdhw7b3aBX5QtuaVEEUhp8UcwjSVjiSusOxC9HT0a2kkMe2F27QCOwoEOS91
JvmRv2IqwgF0ObY4Ymk7npx/pDpWnhJj3f3/PdD/uLlt+hDNnr74tFRmaIizRmfN
kh0jlJLgN3pAkRJUJNPowKmgMe7rKSEbmHQiJGLAd2eaA4lwhT789fWPfKfKhr1t
A739PzM3nKj6wZlQGOTwilQDy9xgoQgvanu8zvkcJzbdblD8Q6Gq4NrNNwGVQntJ
jpZvksNP6YvTlQwKgT3lFELWhEUFJXhKv3QSLBhal4lvQwUxRSXszLnBjhLpQ25K
B0dXXW/VM1UWWMb+4klo+NP6E7KyeorN4xtgknQBrWNLMUz45uuHc8bv84cM1ldH
rZM0h3HjBqcDjGJr8OUnNxUNrqVbbVXjMBqc49UWR58gJ4Bj+WTVM3pizxRBodzT
WZuv/4qtEn/xbOSiyJzobdlIZORMpmnACIrDaZMfEHjoTZWqvfONX+uZw1lzzkZz
Xtvjr7EKOcN6yc25QT+053Yhi/s4BpeXborJkZAxBrFgMy85+5JeGTGAbnB4NvoE
UaMAo1KiS7+nM3JUJapbucbnAe2ZvHfrBTk3pYs23lH8UPm5/bsr8Oy55UU4JAQ4
pt+IwltVHj2IToDJ4BGGeSoNtzcsyamGbSljpMbBuHlwlfFlCZa6fEe9IyQuvnYY
OAHAxATBNFB6pVNUEzPpBGXuS6rOM/JSDeY6o9NEUj62xO+Sdy0+e9N2exz0Nd5l
GXaNbv2mnJBG5I1cmI0yBYNpN85ylFlUgr3rdkzGyF5UtMltnDsw+GG5L4PAI9si
OdYnL4Y5ASsBUqYkGp24thVMCBQuZx1PmWsaPh80T8tu0qAW3nzWNMjniFmeX4Ww
M7B2VB1r0Qi5RbKxEqdyPl+GQ6ny6kBhzGifgitwsEhh2UbxhN4IrOdYDOZH+8z6
qtm0KBFxE8pCM53zOa26Vbu4XtUXM9dwOdtj2pXd81SacRyCrgraK72Pj6X7QIbx
t4OJgjNiminGwRM5ioqvFhoSGOWf3PSSs1F46cSFHrx2Sy1Zw8TdxVF9wpRiVzD/
1SQduPz/+mWZlAizljarNHF7jecU0zsHrUVwteCLpgdi4mnxbtrL7vjxiQ29jblH
Hj5jG6u0kB9Oi8OZP2fOyM6tixo3Z5hy9CcBSYGfqYv50+ZTQr2F6YEuhXKwBayR
eZlxmgy/XbwCFgIeQQnB2YImvTyNJCXMDWyMi1PPYlta+PJBNwaUy43WxuEgxpUG
iOoIea3qwxdUGWCPyVLEzRLe0W0Fs9Fq+rJ1m5Q2/y6l34IRikrzt0N0HO8xAJHz
fsY42g9uqPOv85lvk5Nxw3bqaWUyfQ6OnoPCWimERSGf07F9oGRD0MY6K7Oz1rMn
0JIf4jWef6jyOtmnQOEJpuZ8PlZlZnSEs8zrKvtpa3uCgCWKILvj9+k2cD42Sg9g
GVcgXaIm4b1nfK9h3CZrSbvI52t8Uv6yVHeFfjmxbG44yfozExB1nG/PeEBz7dIm
H1noaouaXadupktgHWjywexHe0lUROuQaktezTDyfsqBUJKZ2qeiyez6IWxOK7tu
m4cHcZq4UlG22tcR/SeGpBC3s2De90MaCROZOKMV+JkLfZ+VERhbj44AJIa5/CwU
Od11N6F7hDXRqvgaR0QqjONUOc7lcQtjhVS8ebDRy6EVwugR0kB+FgZDvzDB9cDq
84+GZp7V6dyQqX9KXt4W5MgvFJDUPI/+d+qV0tXJy66u2N86xbkwoZeEo/yk2p2F
AstBPECPYuGoYL+Gz9EL5EpxwQeLkWdzzJl6ePk310mLQwmpdjaH0iAhVQ8Uv1Pg
7Dzw5qtVGNkhGX0FAcgBIO6mPa1A2hXkCpJoRBUzpc6k0P6JaryDBBFeoj4aHLxL
H6iR2cXtORCAfYf0PEe/gOAX/EzjyU+eUg1ny6NXrA5lgCZTCKlDmO2I97FQw0RZ
EI4zVD5Pr3D70VOIa/n+bxZIJNu8rDVcwyiVizfHEUSOsriaO4If/t0zSC5jzvW3
cHP7UTamTRgAO3hn4UtlVdfEWxJsGe7ZLJ8435B504NDyJkSSnp+MLphHFMBjJ+f
Om6PgXOqxOQXX40sijewPGqNu0EBboZZUl7UiLH3ARLDqbkZ+/mge40ach0OTYBd
oFtxOwQjSww4/hpSRijPBmcCDkPId/qWMFIo9/M8fTfOuEtlefGZu9sD69TqIBWP
2Zs8dB4nLhY2IZOegedIjaf4+hVNje7aVvlil4Ba0Cmw7NkRJQttoSlwbhlHvXwH
uYGXLinV2cd/zj8Djbt0vusas/ToFZRnYeE5dTxgrX+O2zV7gk9FIvbuDrNjsc18
CPb+ig8VzBCRCcG0xm7id69IrY7Ea27pW51lNsSFB5Wn8/exEHcRygfeRhVtJqSO
FgPocxQlQCaljoy+AUdUJsOhXOqAkwi/NdyZFT742kOBt6QzKXWGYrNPMbtUq2T5
VXc9UqTztMXYUdnJKYgEjsfuTQugzdhM5BEQwVL5Lrhok43Wrd0odq4LaPIaqXUZ
IAleVM97iVRjHPaSj5DqaPftbdUjBn2RAiqG2jd/sDiLaEB+RY9lQxelq5PoQ2M2
dg1N1RYgflanQeTNU5UyPMRUYQj72oYYblPKCyD0oX8fiChj/2kjkg0qPcUmfcsS
C3Xmr4eXN0K22VJHJFoCoP0sIe0oTJMNE8ub/74R3kJi3nLpM5XXJu2A5cUanMU9
J5tI9WsEn8YEIrAFxpNjJek27J1+4FEQg1sENsRTaO0Jl4LSQxcNIGQJQkDCHhGV
N0Kol0WoWwMvoVrX8x828d3dJK6iOSxA413ExHErz9jWLJZHxc1MokBtJbA8THmo
ja0NE5LH5XuVI6r8k5EAKqjAddTqRRoP0lYRssA0NANJzQK0+V5FMmxMpp0ykxRI
9aqC/TpouKu5qDXeHiocDoIQhNOLMphLu7n0DBZsDnCu1+y4SAxujZEshesvnTjy
J4F4sh49pavZWk0LwkIZlY0X531ThykvEZLKa6oJEWadgjZJQfkfA1PADV9vrg6h
2cGM9rADSIiF6wXypc7FRw4ch/MRlP8OLz8KEDstR7g61bSxYOB3zmMtQ0I6e/GL
2IDGqvYxrxjvVQbdR5PbSg2zfgHtwO7bgSQ4IxXJGA64+pSPe6jKK7gOnPkzxNQx
B++GWjVpqF4jQelJNdDm3qFcPD3V5bgKSabXXBGMjMEmkdQvk+4Tob/YFlyHdtPR
CkGF24S2ATg+IM7PdqWwlDsrohOlpq7iIhvfg/Xsso4JWsX1l4Utp7CZUyJU8JAs
Sb78DX5t1Y14yHLZo5MrwOTaxFwsuQbiKnai9N5xUJn/m/V/+Hj+ZLdYsM+2qLZz
g3Qu2M9MBobt/nqWkjK6fuLZjLV6o82+HoQ31jGrmGn9edj2whwPOj9oEDB+thgv
WrG/TsxXeixqN8Pr6x/laCX/wAz4oReUWp9KT+4l59dy9lFpTm114qbHkzPlOvIQ
7bQDXeew5s/b3+HudLWeiZNQkIlj8OhhQ1exVyDpO/OsE4D/HVkgZ6d7ZIrGdfwJ
dRdH8UGwkb8AfSKZZCQGKh8Ka5Xc7E1H4HaCdv1mcRztr4QpvWLK4BW4ucbYkCPL
FzodIm3lyGbeICHX9UYCyYrJlEkcMXsVowj3ABkjQ7dcH7whs9vfO3im77U7gmXu
sHiccZFM9juoAD1r88PMFAbSXsJLzoPMp2zfkXMnYRU6VgiaOqRPGIV5Mq+eKB89
Q892qpeqvEBtw7cBtp1NkXHCTye/dmH+eKWme+4tI2b0pkd3XEuhu0ObmONO5ULP
676vLKzFiuiUfqVn5xnH8n4mlkMAq9GDQvghZiZUXhUfHL1ycRc0D5E/S4FONdM1
feAHaXxL3TKrI+6ZYp4wn9npRet6GBCd+coiMXBTLBGoLDLnoFgHBG+b/NkCbXdN
Ng0JBM8eHgQLLrVsvlfroKrQWqvscxRgaOESFcQTmgBAN8hOOnu7rG38hVY0JAgN
gRiSmLz+q66qlGJQjRntEgwgMeg3JKr9nYUZ+H74c0f0TeCgehDVty0N6UMDO+64
qcMAa5LF2n1KIOR6gCdqIAZe45J33rp1ub+3+2ZGBD6xTuoLw21Qf7uaB9o3GYG1
jc/7y2+2IvRQ2ALrD2iICJLiBVBqbI8VJnpYi9HvNdygO/8qBB6z54sjJp8Oh/bi
LF18nIQd1lnl2dUZOqcPuQs6TzSwdSCAjvDsbxlyU8cXcknu2gDcmqfxedCbqIFQ
SHIsesvp2uji4Xg+MFKoQ5a3WkE5yQZuMmkF7MpFpyxYTbUVxC7VWQxJjr5LZREE
vV+7BswkE80PmXsrhzPwBczIOMW3kq4LPMCa+YKw1idwUKPOBcHWnDqnOYzFYmWx
ClAeD/ZgLTh+AyPE/HSkBEsIbLYyk/9VNLKeKRqJOB4FL2JWrTUOn73LgJp8UvjL
dZyAIl2EoxvomUafdhmTGTH1lKjE6IfpfqlNSZZvbsWbAyGYDjRsn1g293vRXzKv
zZ1F5DwrV2my3d/ELhKz1zVome17WmAoiq5RUFSiUoYQfnDpv7iciofU/ZKOfQoY
bbI5GODU8VEqN5iADJoLpEPjKggLyyWkMUw4nbsvJ1pZjXTJmpnVc7fV//u7j5Rl
VQtSzt5aQbdNyZRqyIrhYa9qxiv4fW49MTcQJWmvboHlqG8X8Qb6+YD8+5c3rRUW
/EubgOyPcP8bb8OG1GYsrNStyQAcb3cZklq/JVtotG2QBNo1etpLmYzKB/lfus75
RinTxi5MrkwzF0yUOR0vblj0A9n5LhaN3fDmPVxKjqHYqILt/Ixczf22UiTdeV8f
5Kq/tgi8MeusmLYn7QZ3JgZWqNei2Gdbpn9Ku4atkhWSc6cwrI29aq8/wef0hVnB
vaGWNFm3oiJxTIf7PanrZA1wk4J0mV00eTDC87z5Irv31yB6QBJiWjx3qslxjV6u
evLWdKNj70YFxmXLVUPlBJDCbAlr1Yn3kHqqB09BZOAFUASQjTAF+T0fIn6otF4D
zj0RRj2Zr+BmWPkY2CpxtRq7rJ2sOyYAtAk+cAwDc/0DO9NBmbu+K4VUhsK/jaAk
tCLW4seO9y2r8rDLsW7qUDRr2HLvF2ukNVptbpkiUyM5kq133RB0y+KG8cpENI7U
6SLOnmrc/eTiMWbRHvHomdj8r8hv9EKfTQiZSDyIvA3aj2779agGGN9T0lQvdVmQ
Wld7ZpM45TYIqQZE7MbBa9vuHqnxlIYGNjo2sBoRTXGhE6HHLxb47Vbm5pHSS6sR
pd7r0pUYgo8szieL3q/PvqKNGpAvdLWNzNXtyCGkpmqQwDH1rKEXct2+ZimM8HaX
RBUd+k1wtsZcCghC7MEEifoqbHb/kH40AUUxRn9QmzXfrOnf3Oc67L6myM5bX1dz
raBDTtYU4SLVyQHh5iulCAAitGmqSPatxgRF9iP/J4ySx7fSs+BWwA7B8O2QGim5
L0XsGwzmMn6JBTbhLooXgl5uXZCcxvW8OohHp4XzOLPd8C9N6dhEqnFgUZeo5T1d
DR27RUsKDsSNhOf5YuAvKOnDhmPYUSpeYHWBQxHqathN2uucU+Ji/kImMFl25TCL
mllyypecHFVczLM17Y4Zlht5Qa1FsCkHOFBMRmjx+5p26P1BFyeSsbxs6hV1No7K
SfQvXkkUph6195KZPDTfOcn5gz6x7cMXQCPTziTl5IKQ6mtRVHbfYwy1836OoFMq
ii1yj2Yd+3CrbJ45cWUMoEVWCqVtx+rV3i6j2IN/tojsjwYxa64yFVcFR/uzfFf+
SeYnhzJoq7QQk7y4cHwd4zvkmTK3k2gpr+TA63ePAeZgGD0xC/+s2IiEi0DE4c+T
1cYF4y65ZXttYMXbW8m01thTutXFCAXlWC/rqewxtciyBOo66zTP9O9YvhYmSqPS
lKJ+cTbGL0yozSYQioVkpna03RbByCQEbpavBtkkIiUEuFgzv2gl9M+VYjwrt6Vn
UrM6qXfBwHZCIKvMblslUlHq/QI8rLBK3fwWMxJ+QXCC3NJmxi77h0QJL0ytthLw
qWbUA7s1V3ntF2gdT06vhj9znH7BolfQ4TE4BDL4chtXU6PDXX89eTLvxiy+Cyw1
/U4j26kTt5lZroi45qtB8aoG7fSSUV+oeOC4hiTWfYPVACWHEoQ7cnmR7I56G6VV
xLdgvpEPNVZsViLGUQHUHLxdziv6eauUTntmccuqUmpdhShvuaNogdYAS7gxaHTq
FYyKINTlRHCjFzAt3K/z+rKRuVWDZwl8bwUhOquas+qI5IxZXD2+/MHC904XhiQO
IfP6Es4a8FDoVD5FnbIN6n5JuJD/2pm2ss0WCHtkg4opSAyDYPYh9+71p40EkVBb
BaHiw793HXO/HhaTUmVYQa/HN0utdYl/NCSvg5KFv5iSwqMEClOty+pbK8w20SGI
nxy11eYh4GbYPVti3C0euyFEHAiv70xE8S4C7MvSxUpl5IJPoJANZwRNW9p/rxG7
38jevZ+3Ss4Gjo9sx7euTZ3t2uRw8ke/F2JI5Ua4WVIdMEBp5PaZL4ZuK8r2b9AZ
cK4kUOTLbBCgNAzVnbzRsOihBBpZ1VgPs4PDpx8XIGI3+uRurd4vudruS7VUcqOZ
qBUWBFX/lt6QTNWYRG9SSD+5guNp9Qhl6nYISdl3ZrrtVtObrrgtFnSVD3fqxNYJ
yqIi8Hs8zjZkH1ZZIJaeGjVywW+yi7Uut6rWnda1XP5N7EFyP4Kofr5DwgIVcK6i
n/DZ6MWyzPIeHXEQmIAA6QPGaZXWa0hIvehlDwG/5ZoxpyCur6sU9JEv1W1D3pod
zEf4aNWwOGb+QpgCdw13PFcTwzIUTlz6QYtEsy+nfN3L7Da1s2GSNYMRIZb8Xu+9
JizGpxNEC5EzZACC0WRqDkscZEVULji5o2tp3bBLv91mGrVFgD5jxG3gskKsXNJl
mX6vCFNt/H6xLXVvIu+NDd6sIxt1oyP+wLD4zcbHZVDs1agp3je9dYOnaCAeavEy
70w2KvcFEzljQPzgI7Qvv5wE+iamiZZ+XlzdZ/g/ltaCF7rk+obKUnda3AEtOTXr
LVlITHgVblSgW6n2nHy6tjxH03YaRTAQwX1FL3SGmRaI79RM0dg4soKc9bj8nbie
MInJMgjDFrZrVb5KJEvcMKJE/fgYFf8SDk9CJnjdG3hotymxH9vv2D9w1kMXKYrv
MCvDZxQfWAc11ry/UCDs/BT45HER5QYhcmp7E4A+dEUla4PBONYbKs+aXbRDLtld
Hjp5wMT2eHPmR5ktGKvpWlq5VI+QFnugKs24pfxnTslmSkjzk76tpUkZW2u2yJAD
StyekijOSEzMfBMYtyRxFAzVCoZVZC/22j+cEE18SFm/8vai1t1tLh52MCZtJV5h
BReK+U/cTihZrQSQuckftyOgkOujLYfLrYxUy8CnAKx0nDoYJhbtu58F1Mp/vcYq
JMzuzjdFPhsuT0rDfRiDNqUKacnfPIv68DEd9JCbEy20fQE6yTL2LGb5e7BbHZjw
QE6SVOdqAXfbcWAzKbn8q/yMMZlXk0fATbJYj2eYpJ9M8pzy0Ka5/fhfp/CNX0AH
GLSLb593HTDv9mjr4vh6RlFSD6BgtOlqmH4sU7KmTeQkjRHFSYn5ai9iAmRutyPN
+3UTfia0bKJVq1zfwRqmBDaa/zskiYwBcuSp9P0wTNJi9BT/k7px5IG6TzbHqxyl
AKpIEono6d+CJEPlN0PExkfD/xFcIP3ITWusVNqA7AffTR6n7dvMr3KmqnOo9ZI/
kBDJrpYAT5nh/ZUPP4pMuXWIPR2YUFLWHVm9eixhn9jGAShjBq/yAeVsFptfP76E
hKosMjkPwXn72ddWFkpL7hhqP7LlPNsvG5MDzGNmGc9mgNUgjv6ou9og60jbCPWR
KLam2llOZOMyWL8toLqMpUJo0u4kcwfEWboln+W5Z0TrYr2ltUgoEyPYXxKBZW8d
1XLYLWpR4tb1O6h8MASNYipsy91d50ih4DsJHsSIvqiBCxsWONsLkGgXBi+37CQC
IYgMD1lu+EKZHxPHJCmEnWtsisb2D2Vvg9kfESO5Ot/zjAn8M6pfTosuGxjPNSZv
S+fc5IeIyaDOLMsfWKcZKSgGET6O+KvHMSD9w+Z2mZeqLg10vJinL2d6LP9u9USU
o5b0L/dL6FXzNxqtVsTumYJT8jYvy/SPCA3PjOLajjF6OQh17ZJFk1+kEb1YRy67
l3ne/zk0PV6OMScLy8gSxhmKxdKje8sw5aGypFsHWF/w8YOxjUIRQTmFvu2OTMEg
YHdjI/lhQjWmZ55B906f8ceZ2GehFl7DAzC6ZEPl7CCgICRprlz69IkwNAwYWp0c
YVqgPSCpmIrWgkTfN4It6uwQz53WRORRCZaS0r26OPGXrE9l4du5kM7Mgx/oVMqc
VpX8iaNy56mWxJd8e863a1o95g3lP1uy1sVkjAslAtr3R6/87v7UHY4QqjjwDYnR
2hRqw3T6vDwKO1u/2eDKIGBth9gvDIXw8A/aVOO/6tuDySslBev+mAo7sPFQZ1Eg
DYyn3Rc75GbmgRwokQTUux8AVp5CR1UIKCwsVT3sVB4sa48uiuRs6QytlBcwPCfA
NLQkxCDDSijTYkq+q5nBqCuWfgURvnakZloAAG6wrWItr3uFj8Wr3G90pmjVnmpx
53BSV0Z9Mo3OCca/CVimHA5WEUb0SDvYxX9iSBroDVK4tO0C828CYVbJgLDKFAYn
rQBhFXb5NHtGD8VQ9CmHvrQLBGOOIIYXPB9tIZGsq4PHGsiyuvHAjvD86lFOGsOS
snJYXFT3mCSrAk2qP1gMXZ7csY1pbNk07I9D/uWHfBja1ZG7mG+117NQGBmJEfh4
y/eqklqf7JSrAC0iq2ukO7/ItSQ12h9YppPbVv4Ro7Vj/1pKv2Ef94UVv4QkIQB0
XcPuAchODFx0GWXyiwjIImAti27seHHbH1KEoOYVpU/nbb8qn8jf1S2H368dhe9k
WiRvKn8W0ofbZN8lHllRMsJVHghC+D6BzwtX8iivJo1L6yCdqwH1ln0hirGg3uuU
9yMXr/h0qa9yp9xyl5DsHbSU8iyowcf0m9dRdYQgpcEU5WaU11uN5EwCFI0HMDH6
kSQiQAxxBc1sHQeLrQF1BvjuaBAcOqB/XeaC5wWol2K9f+osuHorJ+7+NLGFCbyN
Tm1IjHiFzawD39CVCcajYBIh2Et+0ZvRitoDwcc0pdGtQHp/WUiVBf/VdOzFKxpu
u8kBykK6B7aFp2NoLbJiXfbqbqaJ+sTI60je8QpbPazUkhaedlEioGKFOV0K9zdb
NFLTQ0tqk7rAvK6dkumPfRDIKxd7NAa9H4sOrbQlR82kIQtPjMUaHfmAZO/40GTq
t7CfYzZ5wRUXvDFLtcjvCQTkgdx3cYrPcESsE9qAMWsoCPIfeZesIV4JvUAcQGg3
l44KVI32Gxgri+RYYIEdWdg2sEsxi5staE2rrZJeX7xrC+BAq09FadVeFLeB9Pl2
AgZL1J2mILqjVSS7dL3c4wdD3Prx+249U+5+IiybgO6LjIQi6Gf2szynSsszSFXT
xKCdwaqX4I4WNtNtf2u22Q==
`pragma protect end_protected
